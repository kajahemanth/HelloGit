------- Test file -----------
library ieee;
use ieee.std_logic_1164.all;
--------
-- Try to add some sensible code here --
