------- Test file -----------
library ieee;
use ieee.std_logic_1164.all;
--------
-- Try to add some sensible code here --
-- Define Sensible? --
-- Let me say that for now we need to stay calm --
-- Time for a new branch --
-- changes made for merging the main branch --
--- change again just for the depth of the branch--
